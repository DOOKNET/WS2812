module RZ_Control(
	input	clk,
	input	rst_n,
	input	flag,
	output	RGB
);

//----------------------------//
reg 	[23:0]	RGB		//24bit数据，发送顺序：GRB

//----------------------------//




//-----------计数器------------//
always @(posedge clk or negedge rst_n) begin
	if()
end
//----------------------------//




//----------------------------//
//----------------------------//
//----------------------------//
//----------------------------//

endmodule
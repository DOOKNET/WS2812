module RGB_Control(
	input	clk,
	input	rst_n,
	input	symaol,
	output	done_sig,
	output	[23:0]	RGB
);




endmodule

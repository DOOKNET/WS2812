module TOP(
	input	clk,
	input	rst_n,
	output 	RGB
);




endmodule
